
localparam ADD    = 4'h0;
localparam SUB    = 4'h1;
localparam AND    = 4'h2;
localparam OR     = 4'h3;
localparam SHIFT  = 4'h4;
localparam LOAD   = 4'h5;
localparam STORE  = 4'h6;
localparam MOVE   = 4'h7;
localparam JUMP   = 4'h8;
localparam LOADC  = 4'h9;
localparam UNDEF1 = 4'hA;
localparam UNDEF2 = 4'hB;
localparam UNDEF3 = 4'hC;
localparam UNDEF4 = 4'hD;
localparam UNDEF5 = 4'hE;
localparam UNDEF6 = 4'hF;
