
localparam ADD    = 4'h0;
localparam SUB    = 4'h1;
localparam AND    = 4'h2;
localparam OR     = 4'h3;
localparam XOR    = 4'h4;
localparam SHIFT  = 4'h5;
localparam LOAD   = 4'h6;
localparam STORE  = 4'h7;
localparam MOVE   = 4'h8;
localparam JUMP   = 4'h9;
localparam LOADC  = 4'hA;
localparam OUT    = 4'hB;
localparam UNDEF3 = 4'hC;
localparam UNDEF4 = 4'hD;
localparam HALT   = 4'hE;
localparam NOP    = 4'hF;
